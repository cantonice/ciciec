//****************************************Copyright (c)***********************************//
//ԭ�Ӹ����߽�ѧƽ̨��www.yuanzige.com
//����֧�֣�http://www.openedv.com/forum.php
//�Ա����̣�https://zhengdianyuanzi.tmall.com
//��ע΢�Ź���ƽ̨΢�źţ�"����ԭ��"����ѻ�ȡZYNQ & FPGA & STM32 & LINUX���ϡ�
//��Ȩ���У�����ؾ���
//Copyright(C) ����ԭ�� 2023-2033
//All rights reserved
//----------------------------------------------------------------------------------------
// File name:           lcd_rgb_top
// Last modified Date:  2020/05/04 9:19:08
// Last Version:        V1.0
// Descriptions:        lcd��ʾ����ģ��
//                      
//----------------------------------------------------------------------------------------
// Created by:          ����ԭ��
// Created date:        2019/05/04 9:19:08
// Version:             V1.0
// Descriptions:        The original version
//
//----------------------------------------------------------------------------------------
//****************************************************************************************//

module lcd_rgb_top(
    input           sys_clk      ,  //ϵͳʱ��
    input           sys_rst_n,      //��λ�ź�  
    input           sys_init_done, 
    //lcd�ӿ�  
    output          lcd_clk,        //LCD����ʱ��    
    output          lcd_hs,         //LCD ��ͬ���ź�
    output          lcd_vs,         //LCD ��ͬ���ź�
    output          lcd_de,         //LCD ��������ʹ��
    inout   [15:0]  lcd_rgb,        //LCD RGB��ɫ����
    output          lcd_bl,         //LCD ��������ź�
    output          lcd_rst,        //LCD ��λ�ź�
    output          lcd_pclk,       //LCD ����ʱ��
    output  [15:0]  lcd_id,         //LCD��ID  
    output          out_vsync,      //lcd���ź� 
    output  [10:0]  pixel_xpos,     //���ص������
    output  [10:0]  pixel_ypos,     //���ص�������        
    output  [10:0]  h_disp,         //LCD��ˮƽ�ֱ���
    output  [10:0]  v_disp,         //LCD����ֱ�ֱ���         
    input   [15:0]  data_in,        //��������
    output          data_req        //������������
    );

//wire define
wire  [15:0] lcd_data_w  ;          //���ص�����
wire         data_req_w  ;          //�������ص���ɫ�������� 
wire         data_req_big;          //����640x480�ֱ���lcd���������ź�
wire         data_req_small;        //С��640x480�ֱ���lcd���������ź� 
wire  [15:0] lcd_data;              //ѡ�����������
wire  [15:0] lcd_rgb_o ;            //LCD �����ɫ����
wire  [15:0] lcd_rgb_i ;            //LCD ������ɫ����

//*****************************************************
//**                    main code
//***************************************************** 

//���ִ�С���Ķ����� 
assign data_req = (lcd_id == 16'h4342) ? data_req_small : data_req_big;   
 
//���ִ�С�������� 
assign lcd_data = (lcd_id == 16'h4342) ? data_in : lcd_data_w ;         

//�������ݷ����л�
assign lcd_rgb = lcd_de ?  lcd_rgb_o :  {16{1'bz}};
assign lcd_rgb_i = lcd_rgb;  

//ʱ�ӷ�Ƶģ��    
clk_div u_clk_div(
    .clk                    (sys_clk  ),
    .rst_n                  (sys_rst_n),
    .lcd_id                 (lcd_id   ),
    .lcd_pclk               (lcd_clk  )
    );  

//��LCD IDģ��
rd_id u_rd_id(
    .clk                    (sys_clk  ),
    .rst_n                  (sys_rst_n),
    .lcd_rgb                (lcd_rgb_i),
    .lcd_id                 (lcd_id   )
    );  

//lcd����ģ��
lcd_driver u_lcd_driver(           
    .lcd_pclk       (lcd_clk),    
    .rst_n          (sys_rst_n & sys_init_done), 
    .lcd_id         (lcd_id),   

    .lcd_hs         (lcd_hs),       
    .lcd_vs         (lcd_vs),       
    .lcd_de         (lcd_de),       
    .lcd_rgb        (lcd_rgb_o),
    .lcd_bl         (lcd_bl),
    .lcd_rst        (lcd_rst),
    .lcd_clk        (lcd_pclk),
    
    .pixel_data     (lcd_data), 
    .data_req       (data_req_small),
    .out_vsync      (out_vsync),
    .h_disp         (h_disp),
    .v_disp         (v_disp), 
    .pixel_xpos     (pixel_xpos), 
    .pixel_ypos     (pixel_ypos)
    ); 
 
//lcd��ʾģ�� 
lcd_display u_lcd_display(          
    .lcd_clk        (lcd_clk),    
    .sys_rst_n      (sys_rst_n & sys_init_done),
    .lcd_id         (lcd_id),  
    
    .pixel_xpos     (pixel_xpos),
    .pixel_ypos     (pixel_ypos),
    .h_disp         (h_disp),
    .v_disp         (v_disp), 	
    .cmos_data      (data_in),
    .lcd_data       (lcd_data_w),    
    .data_req       (data_req_big)
    );   
               
endmodule 